module cpu(
    input  wire         clk,
    input  wire         rstn
);

endmodule